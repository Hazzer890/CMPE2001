library verilog;
use verilog.vl_types.all;
entity FDD_Lab2_vlg_vec_tst is
end FDD_Lab2_vlg_vec_tst;
