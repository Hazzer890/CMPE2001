library verilog;
use verilog.vl_types.all;
entity FDD_Lab2_vlg_check_tst is
    port(
        T               : in     vl_logic;
        V               : in     vl_logic;
        W               : in     vl_logic;
        X               : in     vl_logic;
        Y               : in     vl_logic;
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FDD_Lab2_vlg_check_tst;
